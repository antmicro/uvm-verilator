class uvm_reg_block extends uvm_object;

endclass

