class uvm_root extends uvm_component;

endclass
