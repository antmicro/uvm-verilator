class uvm_reg_block extends uvm_object;
   uvm_object_string_pool #(string) hdl_paths_pool;
endclass
